library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity EX_manager is
end EX_manager;

architecture behavioral of EX_manager is

begin

end architecture ; -- behavioral