library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity ME_manager is
end ME_manager;

architecture behavioral of ME_manager is

begin

end architecture ; -- behavioral