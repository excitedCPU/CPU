library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity ram is
end ram;

architecture behavioral of ram is

begin

end architecture ; -- behavioral