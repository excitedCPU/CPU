library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity EX_ME is
end EX_ME;

architecture behavioral of EX_ME is

begin

end architecture ; -- behavioral