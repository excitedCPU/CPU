library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity mux_writeRamData is
end mux_writeRamData;

architecture behavioral of mux_writeRamData is

begin

end architecture ; -- behavioral