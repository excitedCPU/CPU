library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity EX_WB is
end EX_WB;

architecture behavioral of EX_WB is

begin

end architecture ; -- behavioral