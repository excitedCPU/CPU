library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity alu is
end alu;

architecture behavioral of alu is

begin

end architecture ; -- behavioral