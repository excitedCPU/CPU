library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity SP is
end SP;

architecture behavioral of SP is

begin

end architecture ; -- behavioral