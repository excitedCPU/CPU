library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity mux_PC is
end mux_PC;

architecture behavioral of mux_PC is

begin

end architecture ; -- behavioral