library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity WB_manager is
end WB_manager;

architecture behavioral of WB_manager is

begin

end architecture ; -- behavioral