library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity mux_ALUsrc1 is
end mux_ALUsrc1;

architecture behavioral of mux_ALUsrc1 is

begin

end architecture ; -- behavioral