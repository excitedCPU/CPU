library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity mux_wbData is
end mux_wbData;

architecture behavioral of mux_wbData is

begin

end architecture ; -- behavioral