library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity IF_ID is
end IF_ID;

architecture behavioral of IF_ID is

begin

end architecture ; -- behavioral