library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity immediateExpansion is
end immediateExpansion;

architecture behavioral of immediateExpansion is

begin

end architecture ; -- behavioral