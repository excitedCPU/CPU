library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity ID_EX is
end ID_EX;

architecture behavioral of ID_EX is

begin

end architecture ; -- behavioral