library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity branchControl is
end branchControl;

architecture behavioral of branchControl is

begin

end architecture ; -- behavioral