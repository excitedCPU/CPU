library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity riskCheck is
end riskCheck;

architecture behavioral of riskCheck is

begin

end architecture ; -- behavioral