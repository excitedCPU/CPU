library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity commonRegister is
end commonRegister;

architecture behavioral of commonRegister is

begin

end architecture ; -- behavioral