library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity IF_manager is
end IF_manager;

architecture behavioral of IF_manager is

begin

end architecture ; -- behavioral