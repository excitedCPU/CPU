library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity instructionRegister is
end instructionRegister;

architecture behavioral of instructionRegister is

begin

end architecture ; -- behavioral