library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity T is
end T;

architecture behavioral of T is

begin

end architecture ; -- behavioral