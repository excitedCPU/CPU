library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity controlUnit is
end controlUnit;

architecture behavioral of controlUnit is

begin

end architecture ; -- behavioral