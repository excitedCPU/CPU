library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity ID_manager is
end ID_manager;

architecture behavioral of ID_manager is

begin

end architecture ; -- behavioral