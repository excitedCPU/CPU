library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity IH is
end IH;

architecture behavioral of IH is

begin

end architecture ; -- behavioral