library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity mux_desRegister is
end mux_desRegister;

architecture behavioral of mux_desRegister is

begin

end architecture ; -- behavioral