library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity mux_ALUsrc2 is
end mux_ALUsrc2;

architecture behavioral of mux_ALUsrc2 is

begin

end architecture ; -- behavioral