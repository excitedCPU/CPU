library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity PC is
end PC;

architecture behavioral of PC is

begin

end architecture ; -- behavioral