library IEEE;
use IEEE.SED_LOGIC_1164.ALL;

entity byPass is
end byPass;

architecture behavioral of byPass is

begin

end architecture ; -- behavioral